`include "uvm_sequence_item"
`include "uvm_sequence"
`include "uvm_sequencer"
`include "uart_tx_config"
`include "uvm_driver"
`include "uvm_monitor"
`include "uvm_agent"
`include "uart_rx_monitor"
`include "uart_rx_agent"
`include "uvm_scoreboard"
`include "uvm_env"
`include "uvm_test"